module counter(out, clk, rst);


endmodule