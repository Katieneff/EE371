module parallel_to_serial(data_out, data_in, counter, load, clk, rst); 
	output reg data_out;
	input clk, rst, load; 
	input [7:0] data_in; 
	input [3:0] counter;
	
	reg [9:0] temp;
	reg [1:0] state;
	
	reg [3:0] count;
	
	parameter OP_NOP = 2'b00;
	parameter OP_COUNTING = 2'b01;

	
	always @(posedge clk) begin
		if (!rst) begin 
	  		temp <= 10'b1000000000; 
			data_out <= 0;
			state <= 0;
			count <= 0;
		end else begin
			case (state)
			
				OP_NOP : begin
					if (load) begin 
						temp[8:1] <= data_in;
						state <= OP_COUNTING;
					end
				end
				
				OP_COUNTING: begin
					data_out <= temp[9];
					temp <= temp << 1;
					count <= count + 1;
					if (count == 9) begin
						state <= OP_NOP;
						count <= 0;
					
					end 
				end
			endcase
		end
	end		
endmodule 
